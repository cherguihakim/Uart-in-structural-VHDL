library verilog;
use verilog.vl_types.all;
entity RTD_vlg_vec_tst is
end RTD_vlg_vec_tst;
