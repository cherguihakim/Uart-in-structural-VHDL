library verilog;
use verilog.vl_types.all;
entity controleur_emetteur_vlg_vec_tst is
end controleur_emetteur_vlg_vec_tst;
