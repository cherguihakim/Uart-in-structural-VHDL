library verilog;
use verilog.vl_types.all;
entity diagram_test_uart_fsm_with_uart_emetteur_vlg_vec_tst is
end diagram_test_uart_fsm_with_uart_emetteur_vlg_vec_tst;
