library verilog;
use verilog.vl_types.all;
entity eight_bit_serial_shift_right_register_vlg_vec_tst is
end eight_bit_serial_shift_right_register_vlg_vec_tst;
