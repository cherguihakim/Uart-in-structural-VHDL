library verilog;
use verilog.vl_types.all;
entity mux_8_a_1_vlg_vec_tst is
end mux_8_a_1_vlg_vec_tst;
