library verilog;
use verilog.vl_types.all;
entity UART_FSM_vlg_vec_tst is
end UART_FSM_vlg_vec_tst;
