library verilog;
use verilog.vl_types.all;
entity baud_generator_vlg_vec_tst is
end baud_generator_vlg_vec_tst;
