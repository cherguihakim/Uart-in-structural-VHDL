library verilog;
use verilog.vl_types.all;
entity UART_EMETTEUR_vlg_vec_tst is
end UART_EMETTEUR_vlg_vec_tst;
