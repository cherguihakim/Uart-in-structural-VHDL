library verilog;
use verilog.vl_types.all;
entity diagram_test_uart_fsm_with_uart_emetteur_vlg_check_tst is
    port(
        o_TxD           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end diagram_test_uart_fsm_with_uart_emetteur_vlg_check_tst;
