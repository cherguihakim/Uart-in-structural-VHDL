library verilog;
use verilog.vl_types.all;
entity RDTD_vlg_vec_tst is
end RDTD_vlg_vec_tst;
